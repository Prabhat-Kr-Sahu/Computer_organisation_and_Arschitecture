// pc.v neutralized
// The active `pc_update` module implementation is in `pc_update.v`.
// This file intentionally left blank to avoid duplicate module definitions
// that cause elaboration errors when the simulator/synthesis tool finds
// multiple modules with the same name.
